library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


Entity FirstPipe is
port (
	Clk,Rst:in std_logic;
	PC_Sel:in std_logic_vector(1 downto 0);
	PC_Plus,Jump_Rdst,RET_RTI,Call_Dst: in std_logic_vector(15 downto 0);
	PC_PlusNew,Instruction: out std_logic_vector(15 downto 0)
);
end entity ;

architecture FirstPipeArch of FirstPipe is

component my_adder is 
port( 
	a: in std_logic_vector(15 downto 0);
	s : out std_logic_vector(15 downto 0));
end component;

component mux_4to1 is
  Port ( SEL : in  STD_LOGIC_VECTOR (1 downto 0);     -- select input
           A,B,C,D   : in  STD_LOGIC_VECTOR (15 downto 0);     -- inputs
           X   : out STD_LOGIC_VECTOR (15 downto 0));-- output
end component;

component syncram is
Generic ( n : integer := 10);
port (
clk : in std_logic;
we : in std_logic;
PC : in std_logic_vector(15 downto 0);
--datain : in std_logic_vector(15 downto 0);
Instruction : out std_logic_vector(15 downto 0) );
end component;

component my_nDFF  is
port( Clk,Rst : in std_logic;
d : in std_logic_vector(15 downto 0);
q : out std_logic_vector(15 downto 0));
end component;

signal Mux_Out,PC_RegOut: std_logic_vector(15 downto 0);

begin
Mux: mux_4to1 port map(PC_Sel,PC_Plus,Jump_Rdst,RET_RTI,Call_Dst,Mux_Out);
PC:  my_nDFF  port map(Clk,Rst,Mux_Out,PC_RegOut);
Adder: my_adder port map(PC_RegOut,PC_PlusNew);
Instruction_mem : syncram generic map(n=>10) port map(Clk,'0',PC_RegOut,Instruction);



end architecture;