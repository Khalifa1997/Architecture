library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mux_4to1 is
    Port ( SEL : in  STD_LOGIC_VECTOR (1 downto 0);     -- select input
           A,B,C,D   : in  STD_LOGIC_VECTOR (15 downto 0);     -- inputs
           X   : out STD_LOGIC_VECTOR (15 downto 0));-- output
end mux_4to1;

architecture Behavioral of mux_4to1 is
begin
    X <= A when SEL = "00" else
         B when SEL = "01" else
         C when SEL = "10" else
         D ;
end Behavioral;
